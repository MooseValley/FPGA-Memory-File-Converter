BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000500010000010001000F00020100010000000500010001000004040",
      INIT_05 => X"1000100010100000501000001000000010001000F0000010100000F000000010",
      INIT_06 => X"1000100010001000101000004000008000500080000080004000008000008000",
      INIT_07 => X"0010100000100000100000000000101000001000001000000000501010000010",
      INIT_08 => X"1000401010100000101000500010001000100000002000100010000040001000",
      INIT_09 => X"1001010101010101000100000400010000000100040001000100010000010100",
      INIT_0A => X"0001010001000100000100000201001010101010101000000010000010100010",
      INIT_0B => X"0010000010000000004000100010000000000010000040000000000000001000",
      INIT_0C => X"0000500000000040000000000040000000505000100000100000400010001010",
      INIT_0D => X"00100000100040001010001010000000100040001000000000000000000000F0",
      INIT_0E => X"000000000010F000000000F00010000010005020100000000010000010001000",
      INIT_0F => X"5000100000000010000010001000400000000000000000005050000001000000",
      INIT_10 => X"0000000000040000000F01000000000000000000000000010000000004000000",
      INIT_11 => X"0000000000000100000100000007010000000100000000050000000004040000",
      INIT_12 => X"0000040001000001000000000000010000010101000000040300000010100000",
      INIT_13 => X"000010001000F01000001010000010000000F010001000001000100010000010",
      INIT_14 => X"0010001000101001010001000400000000000004000100001000100000100040",
      INIT_15 => X"0000000000005000100010000000000010000000000000000000201000001000",
      INIT_16 => X"0000000010007000000070001000000000100010001000000000501000000010",
      INIT_17 => X"0010000000000000000000000000000000000000000000000000001000000060",
      INIT_18 => X"200000100000F000000000001000001000001000000000100101010000000000",
      INIT_19 => X"0000000000000000000100010001010001000101000100050001000000000100",
      INIT_1A => X"0100000000000004000000000000000101000100000100000000000000050000",
      INIT_1B => X"0000000000000400010000010000040000000001000101010100000001000000",
      INIT_1C => X"006000101000100010100010F010000000F00000000000001010F0100000F0F0",
      INIT_1D => X"001010F0001000400000000000000010100000000000F0000000000000005010",
      INIT_1E => X"0010000000400010000000000000000000000010100060001010100000100000",
      INIT_1F => X"1000000000000000100010005000000000004000000000000000000000040000",
      INIT_20 => X"0000000006000000010000000100050001000000010000000000000004050000",
      INIT_21 => X"0000010000060606000100010000000000000000000000040000000000000400",
      INIT_22 => X"0000040000010000000000010000000400000000000000000000000000000000",
      INIT_23 => X"0400000000000000010000000004040000000000000004040100000000050400",
      INIT_24 => X"0000000000020000000100000100000000000400000000010004040100000000",
      INIT_25 => X"01000004000100060100000100000000010F0001010000040400000000010000",
      INIT_26 => X"0100000000010000000000000004000000000000000000000000000000000000",
      INIT_27 => X"0000000000000002010000000100010000000000000004000000000000000100",
      INIT_28 => X"0000000000010000000400000001000101000100000F00010000010000040000",
      INIT_29 => X"0001000000000000040000000001030100000000000000000000000000000000",
      INIT_2A => X"00000001000500000000010000010000000F0000000000010000000000000000",
      INIT_2B => X"0001000000000100010000000400000001000001000001000100000100000000",
      INIT_2C => X"0001000000000000000000000000100000000010004000001000100000000000",
      INIT_2D => X"00000000000000000000100050000000000000F0000000100010000040500000",
      INIT_2E => X"0000000F00000100000001000001000000010001000001010000000100000000",
      INIT_2F => X"00F0000000000000000000001000100000000000001000000000000000100000",
      INIT_30 => X"0010000000000000040000000003070000000000000000000000000000000400",
      INIT_31 => X"0000000400000100000500010000000005000000010000000500000001000000",
      INIT_32 => X"0400000010000000000000000000004000000000000005000000000005010000",
      INIT_33 => X"0100050000010000000400000100040000000000010000000000000000010000",
      INIT_34 => X"0000000000000100000100040000000000000400000000000000000504000000",
      INIT_35 => X"0000000040400000000000000000400010000000001000000000000000000000",
      INIT_36 => X"0000000000000000100040400000000000004000100040401000001000001000",
      INIT_37 => X"0010000000101000001000004000100040001000005000100000100050100040",
      INIT_38 => X"001000000000F000000000000000000000100000100000001010005010100050",
      INIT_39 => X"0010100000100000001000500010000050100040001000401000501000401000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"000000000060008000001030A0A0F000B07030A0A000005000A020A010005050",
      INIT_05 => X"0000A0308080000030A03010000000004020A0A0F00000C08000B0F0F00000C0",
      INIT_06 => X"8000500050005000508000005000A0000090A00020A000009000A00020A00000",
      INIT_07 => X"00A0804020C04010000040100000A0804020F04010000040100080A0804020C0",
      INIT_08 => X"F000E0A080804020C0F0004000B000C00080401000F0000000900000F0000000",
      INIT_09 => X"80060606060606060002010004040F0000040C000D000A040A02000004080C04",
      INIT_0A => X"0208080408020C0A000901000A0D00303030303030F0000040F00000A08040C0",
      INIT_0B => X"40C040408020401000D000C040804010000040C010008000A00000004020F000",
      INIT_0C => X"10002000A0000040A00000100020A00000804000D04020C01000F000C000C0A0",
      INIT_0D => X"00700050F000C000C0C000A080A00050F0003000A00000F0F00040A00020B0F0",
      INIT_0E => X"00A0000050D0F0F00020B0F000F0000020000040A040A00040C00040F050F000",
      INIT_0F => X"0000A040A00040C00040F050F0007000A00040A0000010004040A0040C040100",
      INIT_10 => X"00040A00000C000A000F0A000F00000A000404010000040A0200010007000402",
      INIT_11 => X"0A00040100000F00040B000100020A0404040804040100080A000000030C0A00",
      INIT_12 => X"000007000C0000070004020A00000A000400000A0401000D0F0A0000B0800040",
      INIT_13 => X"2040C00070A0F0B00040C080A000904020A0F0A000D04020C000D040700050F0",
      INIT_14 => X"200000C00080F00A08000D0001000A0004010001000C0040C000A04050F00010",
      INIT_15 => X"00A0004010000000C000A04040A00050F00000A00000404010004080004080B0",
      INIT_16 => X"0040A000D000C0401000C040D040100000C0408000704040100020C040404080",
      INIT_17 => X"007040401000004040404040100000A00000204010404040100000D040100010",
      INIT_18 => X"90A000A020A0F000A0004020C0A0007000400020A0005080080B0C0A000B000A",
      INIT_19 => X"0000040204020A00050A0008000C0B000800070B00070002000C040A00000D00",
      INIT_1A => X"0000040A0001000B000A00040A00040A08000D00000C04040A00040100020004",
      INIT_1B => X"040A000401000D000A00040700000D000A00040C000B0D0C0700040208050A00",
      INIT_1C => X"00E000C0D000A00070D020A0F08020A000F000A0000040008090F08020A0F0F0",
      INIT_1D => X"008090F040C000D000A00040100000C08020A00040A0F00040A00040100000A0",
      INIT_1E => X"40B00010001000A00020A00020A00040004010F0F0003000B0A0802040A00000",
      INIT_1F => X"7000402040004000F0007000000040A00000500040A00040A0000A00000F000A",
      INIT_20 => X"000401000F0002040D0404040F0002000F040A0008040A00040404000E000004",
      INIT_21 => X"04020D00040D050C000C010F000402010400000A0000000B0A00000402040B04",
      INIT_22 => X"01000100040A020A0004000F04010009000A0000040404000000040402010400",
      INIT_23 => X"0C000A00010000040A00000F000F0C00040A040401000D0508040A0000040C0A",
      INIT_24 => X"0A04040100020A00040A00040700000F010001000A000400000E050A04020A00",
      INIT_25 => X"08040404000F000E0A02040A040A00000D0F000D0904000F0C000404020D0002",
      INIT_26 => X"0C000404010F0004020401040005000A00000F00000A010404040100000A0000",
      INIT_27 => X"000004040401000B0B0004040C000A00040A000501000D000A00040A00040C00",
      INIT_28 => X"040A0004050F00010001000A000D020A080404020A0F000C01000C0100040A00",
      INIT_29 => X"040D0A00040401000504040A000A0F0504020404000A00040402040A0005040A",
      INIT_2A => X"0004020F000200040A000D04020A04040A0F00010000040D0D0D0D0D0D0D040A",
      INIT_2B => X"000A040A00050F040D040100010004040A00020B00000F040000000D00000A00",
      INIT_2C => X"000D000B040A00000B0000A000408000A00000D000E00040C000A040A0004050",
      INIT_2D => X"4040A000002040004050F000200040404020A0F000F000D000F04000103000A0",
      INIT_2E => X"00040A0F04040F0004040F00040F00000005000800000C040000040F0020A000",
      INIT_2F => X"A0F020A00000A000A0000000D000A000A000A00040F050A0000000D000400010",
      INIT_30 => X"40C0E000000401000C000404040306040A000404040A00040404040404000700",
      INIT_31 => X"0401000500040C0B00020A0C0404010008000A050504010004000A0205040100",
      INIT_32 => X"01000A00504010000040A020401000500040A0040100000004040100040F0404",
      INIT_33 => X"0C000300040C0401000900040C000F000A0004040D040100000A0004040D0401",
      INIT_34 => X"00000A0004040D04010800040004040401000500040A0004040100020C00040A",
      INIT_35 => X"00401000E0E00040A0A04040100050008040A00040D00000A0004040100000A0",
      INIT_36 => X"0000F00000A00040F000D01000A00000F000900080005050C00000D00000D000",
      INIT_37 => X"0080100000809000008010001000C0005000C010002000F00000700040000070",
      INIT_38 => X"0000000000A0F00000A0000000A0000000D000000000000000000040C0900050",
      INIT_39 => X"00A0800000D0100000D0005000D0100000A000F000F000405000204000D00000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000400000003070006000F00040600060000000400070000070004050",
      INIT_05 => X"7000700000200000404000702000000070006000F0003070600020F060004070",
      INIT_06 => X"6000300030003000302000004000700000407000007000004000700000700000",
      INIT_07 => X"3070600000700070500000700000706000007000705000007000407060000070",
      INIT_08 => X"0000407060600000700000404040004000700070004040200070000040002000",
      INIT_09 => X"2005050505050505000707000400000000000700020007000700020000070600",
      INIT_0A => X"0006070007000705000707000402004040404040406000000000002070600070",
      INIT_0B => X"0070000070000070002000700070007000200070700040005000000000002000",
      INIT_0C => X"7000400070000040700000700040700000405000200000007000400070006070",
      INIT_0D => X"00600000700040007070007060500000700040007000007060000070000020F0",
      INIT_0E => X"003000000020F060000020F00070002040004040700050000070000070007000",
      INIT_0F => X"4040700050000070000070007000400060000050000070005040700007000700",
      INIT_10 => X"0200070000040007000F02000000000700000007000500070000070004000000",
      INIT_11 => X"0700000700030200000400070007070000000700000700040200000004040200",
      INIT_12 => X"0000040302000002000000040000020000070706000700050507000070600000",
      INIT_13 => X"000070007050F07000007060500060000050F070002000007000200060000060",
      INIT_14 => X"0020007000602007070003000500070000070004000700007000700000000050",
      INIT_15 => X"5070000070005000700070000050000000005020000000007000606000006020",
      INIT_16 => X"0000500060002000700020002000700050700060007000007000207000000060",
      INIT_17 => X"0070000070002000000000007000007000000000700000007000002000700070",
      INIT_18 => X"607000700050F000700000007060002000007000500000700707070700040007",
      INIT_19 => X"0000000000000500000700070007040006000006000000040007000700000200",
      INIT_1A => X"0500000700070004000700000700000706000300000700000500000700040000",
      INIT_1B => X"0005000007000400070000020000040005000007000602050200000007000000",
      INIT_1C => X"006000702000700070200070F060005000F00050000000007020F0600050F0F0",
      INIT_1D => X"007070F0007000400070000070004060600070000050F0000070000070004070",
      INIT_1E => X"0070007000500020000050000070000000007070600060705070600000200000",
      INIT_1F => X"2000000000000000600000005050007000005000007000007000070000040007",
      INIT_20 => X"0000070006020000020000000000050007000700070007000000000004050500",
      INIT_21 => X"0000020000060606000007020000000700000002000000040200000000000400",
      INIT_22 => X"0700050000070007000000070007000500020000000000000000000000070000",
      INIT_23 => X"0400070007000000020000070004040000050000070004040600050000040407",
      INIT_24 => X"0700000700020700000700000200000707000402050F00060005050700000700",
      INIT_25 => X"07000006020000020700000700070000030F0002070000040400000000020000",
      INIT_26 => X"0000000007020000000007000005000700000000000707000000070000020000",
      INIT_27 => X"0000000000070006020000000700070000050000070005000700000700000700",
      INIT_28 => X"0007000000060007000400070002000706000700050F00070700070700040700",
      INIT_29 => X"000205000000070004000007000700020000000000050F000000000500000007",
      INIT_2A => X"00000000000400000700020000070000050F0007000500030303030303030007",
      INIT_2B => X"0007000500000700020007000400000002000007000007000500000300040700",
      INIT_2C => X"0002000700070000020000700000200070000030004000007000700070000000",
      INIT_2D => X"00005000000000000000000040500000000050F0007000300000000040400020",
      INIT_2E => X"0000070F00000200000002000002000000020005000007020000000200007000",
      INIT_2F => X"70F0007000007000200000002000700070007000007000200000002000200000",
      INIT_30 => X"0070300000000700040000000005020007000000000700000000000000000400",
      INIT_31 => X"0007000400000705000407070000070004000400040007000400040004000700",
      INIT_32 => X"0400040040007000400070000070004000007000070004050000070004070000",
      INIT_33 => X"0700040000070007000400000700040207000000030007000207000000030007",
      INIT_34 => X"0002070000000300070000040000000007000504000700000007000404000007",
      INIT_35 => X"0000700040400000700000007000400070007000003000207000000070000070",
      INIT_36 => X"0000000000700000700040400020000000005000700050500000003000002000",
      INIT_37 => X"3070700040707000507070005000700050006070004000700000000040000040",
      INIT_38 => X"402000002050F000205000004000000020200000500000507000004070000040",
      INIT_39 => X"0070600020707000402000400020700050000050000000400000400000400000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000F0005000C090009050F000D090009050000040009000509000E040",
      INIT_05 => X"1000900050900000205000909000000090009050F000E040100090F040002040",
      INIT_06 => X"100040004000400040900000B00040000050400000400000D000400000400000",
      INIT_07 => X"C010500000500090C0000090000010500000900090C000009000101050000050",
      INIT_08 => X"500090105050000050500090E01000100090009000D0409000100000D0009000",
      INIT_09 => X"9009090909090909000109000F00050000000D000F0009000100090000090900",
      INIT_0A => X"000909000900050D000909000D0900D0D0D0D0D0D0500000005000A010500090",
      INIT_0B => X"005000009000009000F000900090009000F00050900030005000000000009000",
      INIT_0C => X"9000500040000010400000900090400000505000D00000509000D00090009010",
      INIT_0D => X"00000000C00090005050001050D00000C00010000000005050000040000090F0",
      INIT_0E => X"00C0000000C0F040000090F000D000F08000E0B010005000009000009000D000",
      INIT_0F => X"E0B010005000009000009000D0009000D0000050000090008030100005000900",
      INIT_10 => X"03000400000F0004000F09000500000400000009000300090000090009000000",
      INIT_11 => X"09000009000E0900000100090004010000000900000900050900000005010900",
      INIT_12 => X"0000090F09000009000000010000090000010901000900050204000040D00000",
      INIT_13 => X"0000500010D0F04000001090D000100000D0F01000D000005000D00000000010",
      INIT_14 => X"00900050001090090D000C000000090000090008000500009000900000500000",
      INIT_15 => X"30900000900090009000400000D0000050002090000000009000F01000009090",
      INIT_16 => X"0000D000100020009000200050009000209000D0009000009000E090000000D0",
      INIT_17 => X"009000009000E00000000000900000400000000090000000900000D000900000",
      INIT_18 => X"5040009000C0F0009000000090D0009000009000D00000C00901090400010004",
      INIT_19 => X"0000000000000D000001000D0009010001000501000500010009000400000C00",
      INIT_1A => X"0C0000040009000F000900000900000105000C00000500000D000009000F0000",
      INIT_1B => X"000D00000900010004000009000001000500000900010D0D090000000C000500",
      INIT_1C => X"00900050C000400010D00040F09000C000F000C000000000D090F04000C0F0F0",
      INIT_1D => X"00D0C0F00050001000900000900080D05000900000C0F0000090000090001090",
      INIT_1E => X"004000900040009000001000009000000000901080003040D010500000900000",
      INIT_1F => X"9000000000000000D00050008040004000005000009000004000040000020009",
      INIT_20 => X"0000090002020000050000000500020009000400090009000000000009020400",
      INIT_21 => X"00000C00000F0C0E0005090900000009000000090000000F0900000000000F00",
      INIT_22 => X"0900060000040009000000090009000500090000000000000000000000090000",
      INIT_23 => X"0C000400090000000900000400030900000D000009000F0C09000D0000090109",
      INIT_24 => X"09000009000C0900000400000900000909000309040F00010005050900000400",
      INIT_25 => X"090000050005000C04000009000400000C0F000D0400000309000000000C0000",
      INIT_26 => X"0500000009090000000009000006000400000500000909000000090000090000",
      INIT_27 => X"000000000009000D0900000009000400000D0000090005000400000900000900",
      INIT_28 => X"0009000000000009000E0009000D0001050009000D0F00050900050900090900",
      INIT_29 => X"000505000000090005000001000400090000000000050F000000000D00000009",
      INIT_2A => X"00000005000F000009000D00000900000D0F0009000300040404040404040001",
      INIT_2B => X"0009000D000009000D0009000500000009000004000009000C00000C000B0400",
      INIT_2C => X"000D0001000400000900004000009000400000C0005000009000400010000000",
      INIT_2D => X"0000D0000000000000005000F04000000000D0F0004000C00050000090F00090",
      INIT_2E => X"0000090F00000900000009000008000000090005000005090000000900009000",
      INIT_2F => X"90F000900000900090000000C000100010009000009000800000009000800000",
      INIT_30 => X"00508000000009000F0000000000000009000000000900000000000000000500",
      INIT_31 => X"000900080000050C000F09090000090005000100010009000E00010001000900",
      INIT_32 => X"0700010010009000600090000090008000009000090005040000090006090000",
      INIT_33 => X"05000C00000500090008000005000202090000000D00090002090000000D0009",
      INIT_34 => X"0002090000000D000905000F0000000009000205000900000009000102000009",
      INIT_35 => X"00009000F0100000904000009000F0009000400000C000809000000090000040",
      INIT_36 => X"0000500000900000C000D0900090000050008000C0008040500000C00000C000",
      INIT_37 => X"E050900000500000205090007000500060009090004000C000005000F0500050",
      INIT_38 => X"50900000D0C0F000B0C00000C050000010D00000C0000020105000F010500040",
      INIT_39 => X"0010500010009000004000F00050900050500020005000E05000F05000F05000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"00000000004050E00030E00040E0F00050E00040E000003000E000E0E0004040",
      INIT_05 => X"0000E000E070000040E000E070000030E00040E0F0004090D00050F010003090",
      INIT_06 => X"D000E000E000E000E05000003000B0000040B00000B000004000B00000F00000",
      INIT_07 => X"50C08000008000E0A00000E00030C0800000E000E0A00000E00040C080000080",
      INIT_08 => X"E00040C080E0000080E000504070007000E000E00050407000D0000020007000",
      INIT_09 => X"E006060606060606000F0E0004000E000200080004040E000E000700000E0E00",
      INIT_0A => X"000C0E000E00080C000E0E0005030030303030303080002000E00040C08000E0",
      INIT_0B => X"00800000E00000E0002040E000E000E000200080E0003050A00000000000E000",
      INIT_0C => X"E0004000B0000050B00000E00050B00000404000E00000E0E0004040E000D0D0",
      INIT_0D => X"00A0000010004000808000C080E0000010005020A00000A0800000B0000070F0",
      INIT_0E => X"00A0000000A0F0A0000070F00080003010005040E000E00000E00000E0008000",
      INIT_0F => X"5040E000E00000E00000E00080004050E00000700000E0004040D00008000E00",
      INIT_10 => X"03000F000004000B000F0D000E00020B0000000E0002000E00000E0005000000",
      INIT_11 => X"0E00000E00020D000007000E00070E0000000E00000E00040D00000004040D00",
      INIT_12 => X"000004050000000B0000000700000E0000000E0E000E0004040B000090D00000",
      INIT_13 => X"00008000D0E0F0B00000D0C0C000A00000C0F0D000E000008000E000A00000A0",
      INIT_14 => X"0070008000F0E00E0F00010005040E00000E000405080000E000E00000E00050",
      INIT_15 => X"40E00000E0005000E000B00000E00000E00040E000000000E00060A00000C050",
      INIT_16 => X"0000700090002000E0002000C000E00020E0000000E00000E00050E000000000",
      INIT_17 => X"00E00000E000500000000000E00020B000000000E0000000E00030E000E00020",
      INIT_18 => X"70F000E000A0F000E0000000E0D000700000E000E00000A00E0D0E0B0007000B",
      INIT_19 => X"0000000000000E00000E000A000E070000000E00000E0005040E000B00000A00",
      INIT_1A => X"0A00000B000E0005040E00000E00000C08000A00000800000E00000E00050000",
      INIT_1B => X"000E00000E0004030B000007000005030E00000E000A0B0D0700000001000E00",
      INIT_1C => X"00600080A000B000D0A000B0F0C000A000F000A000000000C070F01000A0F0F0",
      INIT_1D => X"00C0A0F00080004030E00000E0005080B000E00000A0F00000E00000E00050E0",
      INIT_1E => X"00F000E0006000400000E00000E000000000E0D010006070B0C0800000000000",
      INIT_1F => X"E0000000000000000000E000404000F00000505000E00000F0000F000004050E",
      INIT_20 => X"00000E00060700000C0000000E0004050E0009000E000E000000000002040400",
      INIT_21 => X"00000A0000060606000E0E0E0000000E0000050D000000020D00000000000200",
      INIT_22 => X"0E000400000B000E0000000E000E0005000D00000000000000020000000E0000",
      INIT_23 => X"04050B000E0002000700000F00050505000E00000E0004040D000C000004050E",
      INIT_24 => X"0E00000E00020E00000B00000700000E0E0002040A0F00050003050E00000900",
      INIT_25 => X"0E000007060E00020B00000E000F00000A0F000C0F00000205000000000A0000",
      INIT_26 => X"0E0000000E0E000000000E000004050B00000E00030E0E0000000E00050D0000",
      INIT_27 => X"00030000000E00060E0000000E000B00000E00000E0004000B00000E00000E00",
      INIT_28 => X"000E0000000A000E0003040E000A000C08000E000E0F00080E00080E00020E00",
      INIT_29 => X"000C0E0000000E000500000E000B000400000000000E0F000000000E0000000E",
      INIT_2A => X"0000000E000505000E000E00000E00000E0F000E0002000D0D0D0D0D0D0D000E",
      INIT_2B => X"000E000E00000E000E000E00050000000400000F00000E000A00000100040B00",
      INIT_2C => X"000C000E000F00000D0000F00000D000F000001000500000E000B000E0000000",
      INIT_2D => X"0000A000000000000000E000404000000000A0F000B000A000E00000404000E0",
      INIT_2E => X"00000E0F00000E0000000E00000A000000000000000008050000000E0000E000",
      INIT_2F => X"E0F000E00000E000D0000000A0008000E000E00000E000A0000000D000A06000",
      INIT_30 => X"0080A02000000E0004000000000607000E000000000E00000000000000000404",
      INIT_31 => X"000E00050000080F00040E0E00000E0004000C000E000E0005040C000E000E00",
      INIT_32 => X"04040C00E000E0004000E00000E000404000E0000E00050400000E00040E0000",
      INIT_33 => X"080004000008000E00050400080004050E0000000E000E00020E0000000E000E",
      INIT_34 => X"00020E0000000E000E0E0004000000000E000405000E0000000E00050400000E",
      INIT_35 => X"0000E00040500000E0000000E0004000E000B00000100020E0000000E00050B0",
      INIT_36 => X"0000E00020E000001000404040D00000E000400010004050E000201000401000",
      INIT_37 => X"5080E0005080100030C0E000500080004000D0E0003050100020E00040E00040",
      INIT_38 => X"507000003010F0003010000040E0000020700020A000004000E00050D0E00030",
      INIT_39 => X"00C0800030D0E00030B0004050C0E00040E0004000E00040E00050E00040E000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"6000000000000000000000000000000000000000070707040400070000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000402070100070100070F01050701000700010F00070107070104010",
      INIT_05 => X"200070107000001010701070000010D070100070F0102070200050F07010E070",
      INIT_06 => X"600060006000600070000010F000000010B07000100000105000700010000010",
      INIT_07 => X"50605010106010705000107010C0605010107010705000107010D06070101060",
      INIT_08 => X"7010D060707010106070107090200020007010701050F07000601010F0007000",
      INIT_09 => X"7005050505050502000607010D0107010F0100010D0407010701070001070701",
      INIT_0A => X"0105070107010607000707010504004040404040400010A0107010D060501070",
      INIT_0B => X"106010107010107010A040701070107010A010607010E0202000000010107000",
      INIT_0C => X"7010800000001000200000702040000020003000701020707020305070202030",
      INIT_0D => X"00500020702060006060206070700020702000402000007070201070002030F0",
      INIT_0E => X"205000002050F070002030F02000204070205030701070002070201070200020",
      INIT_0F => X"5030701070002070201070200020404070001020000070205010600106020702",
      INIT_10 => X"0C02000002080002000F03000702030700020207020302070202070203000102",
      INIT_11 => X"07000207020302000202000702030701020207020207020803000002040D0300",
      INIT_12 => X"00020404050000070001020200000700010607070107020E0507000070200010",
      INIT_13 => X"202060006070F02000106040700070103070F020007020306000701050002070",
      INIT_14 => X"3070006030707007060007020305070001070303030600107030701030703030",
      INIT_15 => X"5070003070304000703070101070003070303070000010107030407000206070",
      INIT_16 => X"00207000703040307030E03060307030E0702050007030307030507020202050",
      INIT_17 => X"0070303070305020202030307030E02000003030702030307030F07030703080",
      INIT_18 => X"306000703070F000700010307020007000107030700030600706070600020002",
      INIT_19 => X"0000010301030700030703020007020005000705000703000507020500000700",
      INIT_1A => X"05000305000703040E0700030700010606000200000602020700020703070003",
      INIT_1B => X"0207000207030E0E020002000003030F07000207030706020700010307030700",
      INIT_1C => X"306000607000700060704020F050407000F04070000030407070F0704050F0F0",
      INIT_1D => X"407050F0306040E0F07000407040E070504070001070F0001070001070404070",
      INIT_1E => X"1020007040B00070004070004070004040407060704010007060504010500000",
      INIT_1F => X"7000104040404040500070405030407000401090207000407000000004010407",
      INIT_20 => X"0002070401040403060304030704050207030700070307000103040404050504",
      INIT_21 => X"010405000403090F000707070002040704040B030400040E0204000104030003",
      INIT_22 => X"0704050003070407000204070407040100030000040404040407030404070404",
      INIT_23 => X"0104050007040C0202000000040B000D040700040704030902040000040C0207",
      INIT_24 => X"070404070404070003020002020000070705080C040F0004050F010704050700",
      INIT_25 => X"07030302060705040705050703060000050F0007000405040000040105050005",
      INIT_26 => X"070505040707000205050704050F0402000007050B070704040507050D030500",
      INIT_27 => X"050A030505070504070003030705020003070005070504000700020700010705",
      INIT_28 => X"0307000505070007050E05070007050607030705070F050607050607050E0700",
      INIT_29 => X"020607000303070503040307000600070005030305070F050105050700050107",
      INIT_2A => X"00010507050703030700070105070305070F0507050E02030303030303030207",
      INIT_2B => X"00070307000507020703070502000201070005020005070205000007050F0700",
      INIT_2C => X"0002000702020000030000700040300060000070503000307060702070002060",
      INIT_2D => X"20302000006030603060706060503040106020F0006000700070406040E00070",
      INIT_2E => X"0001070F01010700010107000105000000070002000006050000010700607000",
      INIT_2F => X"70F0607000607000300000007000500070007000107060700000002000705000",
      INIT_30 => X"106020000101070603000603030501020700020202070002020203030406020E",
      INIT_31 => X"020706040006060006060707040607060E00040007040706050C040007040706",
      INIT_32 => X"010E040070407060906070004070601040607004070602010606070601070606",
      INIT_33 => X"0606050006060607060705060606010407040502070507060407030502070507",
      INIT_34 => X"060E070305020705070707030003050507070304070707050407070601000707",
      INIT_35 => X"0040707030400070700040407070400070507000307070E0700030307070C020",
      INIT_36 => X"0000707080700030707090405020000070705000707050507070107070007070",
      INIT_37 => X"2060707020607070E060707030006070F00060707020007070B07070E07070E0",
      INIT_38 => X"400000701070F0701070007020700070B03070D0500070F06070702060707020",
      INIT_39 => X"0060007020607070200070304060707040707040007070107070807070307000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"80000000000000000000000000000000000008000C0C0C0A0D000C0000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000004090000090005090F00000901050900000005090109090100040",
      INIT_05 => X"9000902090500010009020905000200090205090F020001090F0000090300010",
      INIT_06 => X"80F080F080F080F01050F0300050500040009000405000400050900050500050",
      INIT_07 => X"0090100060500090D0000090500090100070900090D000009060009090607050",
      INIT_08 => X"9070009010906080509070004090009000905090800040500010909000401000",
      INIT_09 => X"9009090909090909000109090009090A0009050A00040900090B010001090900",
      INIT_0A => X"0B0D0909090C05050009090B000D00D0D0D0D0D0D050C000C090D00090100090",
      INIT_0B => X"205020C090E01090D0004090D090B090E000E05090E000408070702080F09050",
      INIT_0C => X"90F000405020F00090205090000050200000404090101090900000509020D0C0",
      INIT_0D => X"00D000109010004050502090409000209020004090002000104030902030D0F0",
      INIT_0E => X"40D00000304000402040D0F04050200090400040903090104090503090505040",
      INIT_0F => X"0040903090F04090603090605050004090006090003090600050100905060907",
      INIT_10 => X"0000050207000409020F0D02090800090207080908000809090909090004000A",
      INIT_11 => X"0902080909000D02000900090A000902070909090A090A000C01020B00040C00",
      INIT_12 => X"020B00040C03000900060D09000009000601090905090C000400020010C02020",
      INIT_13 => X"E0B040001090F09020201010500010100090F0C02090C000402090D0D000F010",
      INIT_14 => X"0090005000D090090002090D0004090205090000050400709010905010901000",
      INIT_15 => X"4090201090100040902090F05090002090200090000050509030000030501090",
      INIT_16 => X"F04010000030003090400030502090400090A0C000902020904000907090A0C0",
      INIT_17 => X"009020209050007090A00020906000902000706090A000209060009060907000",
      INIT_18 => X"70D02090B040F0209020209090D0209000009090900080800901090D02090009",
      INIT_19 => X"0202020A000A090009090A09000909000C00090C000907000509000C02020402",
      INIT_1A => X"0D00080C02090B000409020B090107090803090300050100090003090C00040B",
      INIT_1B => X"00090003090D000409010405000E0004090104090F01010D0900010F090F0900",
      INIT_1C => X"E000605040200000109010903010109000F010400020F0105010F09020D0F0F0",
      INIT_1D => X"0050D0F0E04000004090200090200010103090005090F0205090005090200090",
      INIT_1E => X"5090009030005090005090005090203050209010904000609090106040C02000",
      INIT_1F => X"9050506030604050C0009050004050C02060005000905050C020050207000509",
      INIT_20 => X"0201090700070803050208030908000409000103090209030503080800050502",
      INIT_21 => X"010A05040800070207090909030D0B090909080C0A020B000D0A02020C040003",
      INIT_22 => X"090B00040C090C0902010C090B090C00050D08020B070C0D0D000C020D09090D",
      INIT_23 => X"00040C02090E0000090002050E0804040D09000E090E00050D0E05000F080409",
      INIT_24 => X"090E0E090F0009020D090F040900020909000004010F00000100040902020103",
      INIT_25 => X"0902040006090100090301090E0802020C0F0205050902000404020104050804",
      INIT_26 => X"0904010E0909030D0400090903000509020209040809090E0B050905000C0302",
      INIT_27 => X"05000C02050906000900050009070900050900060906000501020B09000A0908",
      INIT_28 => X"03090006080402090700040902090909090E0909090F09050908050908000903",
      INIT_29 => X"0505090102000909000D030902080009000B06000B090F08010B0909000A0409",
      INIT_2A => X"00020A090A000403090209010D090009090F0C090C0000040404040404050009",
      INIT_2B => X"02090709000E09000903090D0004000409010F09000F09000C0002090E000002",
      INIT_2C => X"02090209000902020C02009020C0D02000202090F00040309020907090008010",
      INIT_2D => X"A020900000200020301090100040C020103090F0208020402090902000404090",
      INIT_2E => X"6000090F0000090000000904000004060F010408000005040007000900609030",
      INIT_2F => X"90F0609070609020C06040401040406090009000009070405000304030906000",
      INIT_30 => X"C040804000090903000404030400030B090C070808090208080A02030D080804",
      INIT_31 => X"00090A08040A05050A0809090E0A090A08050100090E090B08040100090E090B",
      INIT_32 => X"0804010090E090C080A09000E090C08040A0900E090D08040C0A090D08090D0A",
      INIT_33 => X"040E08040D050A090E08040C040E0805090801000900090F0809040100090009",
      INIT_34 => X"0F0809040100090009090000040C020509000004010900010E09010004040109",
      INIT_35 => X"00E09010005050109000E0E09020005090109020E09030809020B02090308090",
      INIT_36 => X"20209040809020B09040004050D0802090400050905000409050009050009060",
      INIT_37 => X"0050906000909060005090600050407000501090700040907000907000908000",
      INIT_38 => X"405000800090F080009000800090209000C09000C00090001090900010909000",
      INIT_39 => X"509050A0000090A00050A000405090A00090B0005090B00090B00090B0009000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"D00000000000000000000000000000000000000A010301000200010000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"00000000005010E01020E090E0E0F05030E000E0E010C04000E080E0E0307070",
      INIT_05 => X"7010E010E0E010A030E080E0E0104010E0F0E0E0F0B0209050F0E000E0202090",
      INIT_06 => X"A0F0A0F0A0F0A0F090E0F0A04090E0208030E020E0E030D04040E01060E01040",
      INIT_07 => X"20D0E06040F060E0E01060E0C010D0E06010E060E0E01060E09030D0E0A0C0E0",
      INIT_08 => X"E06030D0D0E0A050E0E0E0608070107010E0D0E07060D0C01080E0104040D010",
      INIT_09 => X"E00606060606060401090E08030A0E09010A0E0D050F0E060E0B0E010C0E0E06",
      INIT_0A => X"0F0E0E030E070008010E0E010303003030303030C0E09010A0E04020D0E060E0",
      INIT_0B => X"50E050A0E040C0E08050F0E090E030E0602080F0E0E05010A0F0F00090D0E0F0",
      INIT_0C => X"E0304050E070F030707000E04030E040A0805050E05050E0E0E05060E00080A0",
      INIT_0D => X"10E010B0E07040C0C0E0C0D0F0E01080E03050B0D020B0E0E01030E0B0E0E0F0",
      INIT_0E => X"10E0301070E000B0B0A0E0F020E0F020E0C07010E0B0E0F0D0E0A0B0E080E0F0",
      INIT_0F => X"6010E0B0E0F0D0E080B0E060E0D05090E090A0707000E0B0702090030E0D0E05",
      INIT_10 => X"02050E000E040407000F0D000E03010E0507050E0C020D0E08040E03040E0601",
      INIT_11 => X"0E0D050E0A020E000507010E03030E050F040E0C040E0B03010005050709010A",
      INIT_12 => X"050A06090A00010E090A010707010E0A0A050E0E0D0E0007020A050090A040C0",
      INIT_13 => X"5060A01090E0F0E0D0C090708010705070E0F0A050E02030A050E050E01010E0",
      INIT_14 => X"10E010E060F0E00E0A050E0505030E00060E0B05020A0070E0B0E06090E02060",
      INIT_15 => X"30E00040E0E04050E0E0E05060E01090E05020E0A0D06060E01030A000F0D0E0",
      INIT_16 => X"F0D0C010109030A0E05030A08070E09020E0C0A010E00070E0F030E0F04040A0",
      INIT_17 => X"10E00070E09020F04040D070E050104050A04060E0C0D070E0D010E0E0E09070",
      INIT_18 => X"20C0B0E030B0F0B0E000C090E00000E01060E080E010C0100E090E0D0B07010E",
      INIT_19 => X"0B000C05060B0E010B0E0E07010E07010A010E0A010E0E05030E0B0A02030B02",
      INIT_1A => X"0801000F020E0705050E00090E0F0F0D0A000700010E09010E01010E07040409",
      INIT_1B => X"010E01010E0D0505050F0D0E010605050E0F0D0E0D070A000E01050D0E050E00",
      INIT_1C => X"E04040A0F0B0A01090E08050F0E030E010F070B010B000C080D0F0E010E0F0F0",
      INIT_1D => X"9080A0F08010105050E06030E07020D0E0C0E08060E0F00060E08060E0E030E0",
      INIT_1E => X"607010E0E04000E0D030E08010E000F020F0E090E0506050E0D0E080E0A00010",
      INIT_1F => X"E0F0D060F0707090A010E0606050801010C05020B0E00080A0300E020205020E",
      INIT_20 => X"0A010E0E06020C0A0807000A0E05050F0E0D09000E070E0F0602000F0A040209",
      INIT_21 => X"050C0E00070C0000090E0E0E0007010E010D0101000903030E00090C010A0302",
      INIT_22 => X"0E08040C090E0C0E0901050E090E0304040E000404040506000109090F0E010A",
      INIT_23 => X"050F0F070E0101010D01070E07090D050B0E00080E0E07000E080E010707050E",
      INIT_24 => X"0E08080E0E030E020F050F0D0D01070E0E06060C0C0F00010307090E09060900",
      INIT_25 => X"0E070A06050E0A030E060C0E080A07080A0F06080E0108080D050905060E0003",
      INIT_26 => X"0E0505080E0E00070C000E010805020D08060E0E010E0E0804000E0501010B09",
      INIT_27 => X"0D0109090E0E02030E060A0D0E040E090A0E010F0E0804000E05060E080E0E05",
      INIT_28 => X"020E0809010F050E07050D0E060E0B0D0E080E080E0F0A0F0E0E0F0E0A030E00",
      INIT_29 => X"01080E0F070D0E0E030B020E000A000E0006060D0C0E0F0C050C0F0E010E0E0E",
      INIT_2A => X"0D0C0C0E090504020E060E05040E0D0F0E0F0B0E0602050D0D0D0D0D0D0E050E",
      INIT_2B => X"010E0A0E01020E050E020E060404050E0E0A070701000E050A01010E0D020A04",
      INIT_2C => X"030D020E050D04010A0300E020508020A03040E0E0404020E0A0E0F0E070D0F0",
      INIT_2D => X"407050107090D0A020B0E0606070909050B0D0F070A060F080E010D0807050E0",
      INIT_2E => X"50060E0E060D0E030D0D0E030D0A0F0F00000F0A08060B0A03000D0E0020E0F0",
      INIT_2F => X"E0F080E040A0E010A080000080D0A010E0A0E010D0E040D00030009000E0D000",
      INIT_30 => X"A0E0A03000030E0D040400020A07020C0E0D0F0D0D0E0E050D040702020B0509",
      INIT_31 => X"010E01040E030D0E06030E0E08030E0C040408000E080E03050908000E080E0B",
      INIT_32 => X"05090800E080E0302030E00080E0B0501030E0080E02060505080E0A030E0403",
      INIT_33 => X"01000405040E080E06050C0C010D06020E0705010E070E02020E0605010E070E",
      INIT_34 => X"0C020E0A05010E070E0E0504050909000E0F0601010E0D05080E06080905080E",
      INIT_35 => X"0080E0F080304010E0008080E0804030E050E08080E02020E0909070E0B010D0",
      INIT_36 => X"3020E02010E09090E080905040700080E0E04040E0607030E0A010E0E010E010",
      INIT_37 => X"20C0E04020C0E08020C0E0C040001000402090E04050F0E09010E0D030E00060",
      INIT_38 => X"10E0103020E0F08020E010C020E00000201040101010702050E0B03080E0F040",
      INIT_39 => X"00D0E03020F0E08020E0C050E080E0F030E0404000E07030E0B030E0E030E000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

