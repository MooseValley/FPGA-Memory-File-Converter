BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"000000000501001010F0210100050101004410101100510010001010F001100F",
      INIT_01 => X"0001101010101100400805080080400800800110010010000011001001000051",
      INIT_02 => X"1001104111001105010101000201010040101111111101004010001040101010",
      INIT_03 => X"0110011010100100211111111000100110101001000040101000001004000000",
      INIT_04 => X"0100050000400000400055010010040101101001040110110001040100000000",
      INIT_05 => X"00F000001F0000F0100105210000100101050100001001010400000000055001",
      INIT_06 => X"000000004000F100000000000010000400000000010010007100010000500004",
      INIT_07 => X"4000040100100000010011100043001100001010F10011001000F10100101010",
      INIT_08 => X"0101010111101040000004010101001040000005010100000100000000021001",
      INIT_09 => X"0000010700070100001010100005100010100000000000000000000000001000",
      INIT_0A => X"6200100F00000100100100001111000000000000001010110101101050100001",
      INIT_0B => X"0100000040000000110100100000005000000004010010040000101111000100",
      INIT_0C => X"060110101101F1000F00000011F100FF011F010400000001100000F000000051",
      INIT_0D => X"0100040100000000000110601110010010000000101050000040000000000400",
      INIT_0E => X"0000600010001050100010000000450000100666010100000000000400000040",
      INIT_0F => X"0040010000010004000000000000000040000000100004400000004410000540",
      INIT_10 => X"0000020001001000004000010441000010040106100100001F01100440000100",
      INIT_11 => X"1000010000000400000000000000000000000002100010100000004000000010",
      INIT_12 => X"000001000400010110100F010010040001000000400001310000000000000000",
      INIT_13 => X"00010500001001000F0000010000000001000010100040001001001010010000",
      INIT_14 => X"01000000000001000010400101000000000000000105000000F0001010045000",
      INIT_15 => X"00F0010001001000101001100010000F00000000001010000001000000010001",
      INIT_16 => X"0000004000037000000000000000400004001005010000500010005000100040",
      INIT_17 => X"0100000000004000000500000510010500100040010400000100000000100000",
      INIT_18 => X"0001001040000004000000005400000044000000004010000100000000000000",
      INIT_19 => X"0000104400000040104410010010010001100100401040100501001051040100",
      INIT_1A => X"00F0000000000100100011051105011001000105010051040104105104100000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"0000000006080013AAF0B73AA0050A2A105500A388003A31000042AAF00C80BF",
      INIT_01 => X"F00C80505050580050A009A02A0090A02A000A842C41004100A842F41004108A",
      INIT_02 => X"842CF0EA8842CF040B0C08410F000900F00086666666021044F004C0D0A4A200",
      INIT_03 => X"48C4288482CA0910AD333333F004F00A84C4C4482410D0C4841004C1080A0004",
      INIT_04 => X"2F01020A004A00102A00840D42C10F0C0CA0705F0C0CC0A8A05F030A00FF04A0",
      INIT_05 => X"2BF0A005DFF02BF0F002004A4A04C04F5F000A4A04C04F5F070A04A001044A4C",
      INIT_06 => X"41004A00C0A0FA0F00A0441004A20107042A04100F04B0102A444844108A0003",
      INIT_07 => X"CA00070C007042A00A0400A410DFA0B80424C07AFB04C8A0942AFA0D42C0D470",
      INIT_08 => X"5F200C08FA80D010A041010C4C0A45F010A041000C0A44A05F00A00441048048",
      INIT_09 => X"B04A0D0C410C4D4100C480744102C4448074410044444100A00241444100D410",
      INIT_0A => X"19A0A2AF0A042CA070402A0588BCA0B0A004242A05A080CB0807B07020C4A00D",
      INIT_0B => X"0004A010B0A04A04A80D00C44A04102044A0410D0A04700D0A04C0BDC704285A",
      INIT_0C => X"0E0CD0A07D2AF82A0F0A004089F82AFF089F4C0D0A04100C82A04AF04A04100A",
      INIT_0D => X"4B01010A02A02A04041FF030BA824A0070424040F070004A00504A04A0A00F0A",
      INIT_0E => X"0410F024D444F020F4A084A04440E00442D04D5C0C1F0421400A000BA00424B4",
      INIT_0F => X"10104A2A040F41090A00444000442140C0A01004A00F0FC04A4410D584A004CA",
      INIT_10 => X"A44102A04A04700F1010A0400E5A42A084440F0EA24A4A00DF0D940FC0442D02",
      INIT_11 => X"C0441F042414050A00F00A1444100A000044410BB044C0A04A0510D0A04A04C0",
      INIT_12 => X"4A045F01010A0D2A8442AF0C10C104A04DA04410544A0AF542440A04424A054A",
      INIT_13 => X"042F0204A0D42A44AF01004DDDDDDD4A0A4A05F4D4101044A02B00F4000D00A0",
      INIT_14 => X"0D0B4A00B0A0480A00D0E04C0A4A04544A0024045F0204442AF0F0D0F40130A0",
      INIT_15 => X"4AF44F044F04F00050800C4004F2A0AF2A00A0A000D0A0A0A04F5A000D04014C",
      INIT_16 => X"E00410C0444364A0444A0444444070410504CB02AC441080A5541040A2541010",
      INIT_17 => X"A541004A2410504A4100044104F44C0304C410904C0F0A044D4100A044D4100A",
      INIT_18 => X"044D41804044410504A044102C04A410EE04AA44105084A04D00A044100A00F0",
      INIT_19 => X"0A04F0D10A00F0908055C00D00D008100890081010C050C1020F007040070000",
      INIT_1A => X"0AF00A000A000D0000000004C9050A800D100D050D100A0F0F0450240D000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"000000000400037060F0460600040700704570700200440720007060F037602F",
      INIT_01 => X"6047603030303200407004700700407007003760070750070076007075007047",
      INIT_02 => X"6007004766007004440407070442070040202555555507704000007020707020",
      INIT_03 => X"0760067070750770424444446000002760707007007020707070207704050000",
      INIT_04 => X"0207040700470070470045020007040706706007040770765007040700760070",
      INIT_05 => X"02F030002F6002F0702404470500700707044705007007070406005007054707",
      INIT_06 => X"070207004070F200007000705070070400070070320040707700070070420004",
      INIT_07 => X"4200043200200040020077607055707600007075F70076506005F70200702060",
      INIT_08 => X"0602070627703050700704070707000055700705070700500005200007066006",
      INIT_09 => X"2005060207020207057060700702700060700702000007007000070007002070",
      INIT_0A => X"7670705F07000760200705007777704070000005007070740600600040707002",
      INIT_0B => X"0500707040700700760300700500704000500704070020040500706252000700",
      INIT_0C => X"060720707207F6050F05000072F605FF077F070407007046607005F007007047",
      INIT_0D => X"0707050200500700007760675760020020000000600055070050070070700407",
      INIT_0E => X"0070620020000050707070700000455000200666007200070002000420000040",
      INIT_0F => X"7050070700070705020000000000070040707000200704400500704460500447",
      INIT_10 => X"700702700700200770425F060557007070062002700707003F02700440000200",
      INIT_11 => X"0000720000700507000007700070020000000706200070700500705070070070",
      INIT_12 => X"070006070407020760705F07707704700250007040070702000005F000050007",
      INIT_13 => X"00000400702007005F0705033333330707050070207040002007007050030470",
      INIT_14 => X"02070700207002070030400707070000050000000004500005F0703000044020",
      INIT_15 => X"07F0020002002000205007200020707F07007020002070707007020002020007",
      INIT_16 => X"3000704000052070000700000000400704007504770070404040704040407040",
      INIT_17 => X"4407040700704007070450070470070400707040070427000307027000307027",
      INIT_18 => X"0003070040000705407000704400707044007000704070700302700070070000",
      INIT_19 => X"0700704402000050705500030020377047705770507050670407000040044200",
      INIT_1A => X"25F0250040002200500570047004076027704204027050050004004004000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"000000000F050C9095F0D9095004090590E410905900250990009095F0E4109F",
      INIT_01 => X"4024104040404900B04005400400D0400400C1500509C009001500909C009011",
      INIT_02 => X"5005509155005509E10109090D490100D090999999990190F05000D0F0901090",
      INIT_03 => X"09900990905D0990D9DDDDDD500050A1509050090090F0909090F05903050000",
      INIT_04 => X"09090504001400909400550D00590D090910000C09055015D00C010000550040",
      INIT_05 => X"09F0C000CF4009F0D0F80EB1050090090D0EB1050090090D090D005009083105",
      INIT_06 => X"09030400F040F905004000903090090900090090E90010904100090090590005",
      INIT_07 => X"190009F900900010090019109052404D0000501DF40019D0100DF10D0050D000",
      INIT_08 => X"0109050199D0C000900908050909005003900909090400D005029000090F1009",
      INIT_09 => X"900D0102090205090290D090090E9000D090090E00000900400009000900D090",
      INIT_0A => X"054090CF090009D090090D00C91940104000000D0010D091010510501090400C",
      INIT_0B => X"0C004090F0900900150C00500D0090F000D00901040090010500901DD9000C05",
      INIT_0C => X"0905C0401D04F90C0F0C0000D9F40CFF0DCF05010900908D50900CF009009019",
      INIT_0D => X"040904090010090000918034D150090090000000D05084040050090040400209",
      INIT_0E => X"0090220050005020904090900000924000C00FCE059900090009000F900000F0",
      INIT_0F => X"90600409000909050900000000000900C0409000900403900D0090FC90D00919",
      INIT_10 => X"90090C900400900990394F01055900409005050C40090400CF0D400390000C00",
      INIT_11 => X"500099000090060400500990009009000000090D900090400D00905040090090",
      INIT_12 => X"090000090E090D015090DF05905909900550009050010409000005F0000D0009",
      INIT_13 => X"00050F0090D00900DF09030444444401090D0090D090500090040090C00C0B40",
      INIT_14 => X"0D0104009040090400C05009040100000D000000050F40000DF040C05009F090",
      INIT_15 => X"09F0090009008000905005900090909F0900909000C010109009080009080005",
      INIT_16 => X"800090F000000090000900000000500908005C0F99009050101090E010109070",
      INIT_17 => X"1109060900908009090540090690050C00509080050229000D09029000D09029",
      INIT_18 => X"000D0950F00009025090009012009090F100940090F090400C08900090040050",
      INIT_19 => X"0900C0D909005080C084500C00C0E5900500259070506099040C0050F5055900",
      INIT_1A => X"DCF0BC00C5001D00C002150F150401501090040F05905502050E50F50F500000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"00000000045E03E04EF05E04E0030E0EE04400E0E7004E0E7003E04EF049D05F",
      INIT_01 => X"1039D0E0E0E0E50030B004B00B0040B00F005C80080EA00E03C800E0EA00E04C",
      INIT_02 => X"8008E04C8E008E0547070E0E05470D002070E66666660FE040E0208044E0E070",
      INIT_03 => X"0EE00CE0E08C0EE0533333338020E04C80E0800E00E024E0E0E0208E035A0000",
      INIT_04 => X"0E0E040B005B00E05B00440E00EE044E0DD0A001040880C8E001052A00A800B0",
      INIT_05 => X"07F0A000AFA007F08031054E0E00E00E08054E0E00E00E08045E00700E044D08",
      INIT_06 => X"0E030F0040B0FD0E02B000E020E00E05000E00E02D0070E07E000E00E04D0004",
      INIT_07 => X"4D00045000B000700E000EE0E044B09D000080DEFB00DCC0A00CFD0E0080E0A0",
      INIT_08 => X"0A07080FEEF01054E00E04580E0E00E054E00E050E0B00E00E04E0000E06A00C",
      INIT_09 => X"500709020E020C0E02E000E00E05E00000E00E0500000E02B0000E000E03E0E0",
      INIT_0A => X"27F0E0AF0E000ED0700E0E00AEDEB070B000000E00E0A0E7000E00E054E0B00A",
      INIT_0B => X"0A00B0E054E00E00C80A00800E00E05000E00E043B0070053E00E0ABD700010E",
      INIT_0C => X"0608A0B0DA0BFC0A0F0A0000C7F10AFF0CAF08043E00E058B0E00AF00E00E05E",
      INIT_0D => X"0F0E060400E00E0000ED1067BC800000E000000000E0440F00550E00F0F0045E",
      INIT_0E => X"00E06700C000E045E090E0E00000244000A006660EEE000E005D0002D0000020",
      INIT_0F => X"E0400B0E000E0E050D00000002000E0045B0E020700F05550E00E044D0C0045E",
      INIT_10 => X"E00E02E00B00700EE024AF05035E0090E0076E02B00E0F00AF0CF00250000A00",
      INIT_11 => X"E000EE0000E0045B00E03EE000E05D0003000E06E000E0B00E00E040B00E00E0",
      INIT_12 => X"0E000A0E034E0A0C80E0EF08E08E02E00CE000E0500E0B0400000EF0000E000E",
      INIT_13 => X"000E0550E0E00E00EF0E020DDDDDDD0E0E0E00E0E0E05000400F00E0A00104B0",
      INIT_14 => X"0C0E0F00D0F00D0F0010500E0B0E00000A0000000E0440000AF0B0A0E00440E0",
      INIT_15 => X"0EF00E000E00A0000000085000E0E0EF0E00E0D000A080E0E00E0A000D0A6008",
      INIT_16 => X"A200E040000670E0000E00000000440E05008F04EE00E040C0E0E054C0E0E044",
      INIT_17 => X"CE0E040E00E0440E0E05400E04E008040080E05408045E000E0E02E000E0E02E",
      INIT_18 => X"000E0EE040000E0450E000E05400E0E04500E000E040E0B00102E000E05B00E0",
      INIT_19 => X"2E0010444D00E0401045E021041058E058103CE0508040DE035102E04E045700",
      INIT_1A => X"31F031004E002702A0040E05DE030C803DE03B045CE04E040E04E05E04E00000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"600777447427107107F15710701F07177141207170011717001D7107F127205F",
      INIT_01 => X"71E7606060607001F0001B701001507010015651161750171C651171750171D6",
      INIT_02 => X"711671D6771167179202071715F70611F070755555520671D171F101D4717170",
      INIT_03 => X"17711571716707715444444401A171D6517161171171A4717171A1671E220001",
      INIT_04 => X"1707180001020072400203071277235722305027260662677027204200772170",
      INIT_05 => X"23F250025F7023F2024725371702721720253717027217202447012007251616",
      INIT_06 => X"272C20028020F307237022723272272301270272320220723712272272830024",
      INIT_07 => X"D3002445007012200701677172E5707201226067F20164707137F20723607150",
      INIT_08 => X"2737063777607235701733361737137335703734073711703733700117347026",
      INIT_09 => X"70270734373E36373E72507337357222507337352223373E20033723373F7373",
      INIT_0A => X"8360737F07013720701737036767602020013137037320720507507305725007",
      INIT_0B => X"050350734E70370166020062270273703270273EE2020033F702737627013737",
      INIT_0C => X"360670706742F5470F47003477F745FF475F364EF70474E7547017F017017447",
      INIT_0D => X"12074B0704704704447674107654150070144444507453470419270470004147",
      INIT_0E => X"027414436343745273707370134445541450439F0777024744B3404E24014303",
      INIT_0F => X"74503747024747410300444447344744145074C220004B0D4704743924004C27",
      INIT_10 => X"7447447032022007758C4F045F17457073326754755736005F07045400415505",
      INIT_11 => X"7554770255745F420075B7744575D3505A355754703375203705754070270175",
      INIT_12 => X"370557075E57075673757F5675675E702670337534370607053357F515570517",
      INIT_13 => X"01575733707157357F575E233333332707370572737520217052057250075F70",
      INIT_14 => X"02072200307043060075303767270262320063636766534162F060707464E070",
      INIT_15 => X"17F1170117015000702006500176707F67067030007050707017670002075016",
      INIT_16 => X"20117630633512702227022233462E2764066066774676E04074765C4074761E",
      INIT_17 => X"47476967047614674762166761766665066676756661474527576473527576E7",
      INIT_18 => X"352757773035577347775477610774773407704477407570377E703377C20077",
      INIT_19 => X"870377945200775077557717707726772677E6773067F06772077B77E77E4007",
      INIT_1A => X"17F717072707B37D507F67726772060726772073467747740771778773700000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"880CCCADC049009059F0091590005919910490929501092950209259F2019F00",
      INIT_01 => X"93018F8F8F8F15F30550409045040590550509106509D009509107909D009609",
      INIT_02 => X"967597091968597049090959804501990410999999990199099A095A04909B10",
      INIT_03 => X"1990BD999C55099B0DDDDDDD5C0C9D09109252C9E19D049D9B9E0E59E0487728",
      INIT_04 => X"F959F0452F09259005200449119900592DC0D019104552949029204902014392",
      INIT_05 => X"3DF4D00340424DF4520940493914953955404939F49639655049069039605195",
      INIT_06 => X"697005270492FD29809278980899999040A928990D20909A0927999A9A0C12B0",
      INIT_07 => X"4C02B04C30906D90090619959C04021C22EB4019F92211501109FC29C0429DD0",
      INIT_08 => X"F109050D99029D049259005479195191049219104929F5902920900559300351",
      INIT_09 => X"9F41003039403529409AC0922940979AC092295079A02960920769A029609697",
      INIT_0A => X"07D29B4F292299D2900999088919D2909222A0A9099A90990C09C0970590C224",
      INIT_0B => X"2D08C29B0492B9179839305109039C04B09039D0491450E049149F11D901F9F9",
      INIT_0C => X"E0654200191931190F1402F151F92DFF05DFE40049209201139059F259059209",
      INIT_0D => X"59093059059059235291940699164C2095563645C095045C26050955C2527059",
      INIT_0E => X"219707835283980490139293538805521A54807279993DB9998CA2B0DA22C403",
      INIT_0F => X"9B04C9C921C9B9C05D82B7CDD0C2D99D04C29E009025E844D90E9E05DE50F849",
      INIT_10 => X"9EE9F092D9F4902990041F0010492213924069109319E822CF25592044214584",
      INIT_11 => X"941E993D409930592294899EB5950C3250C25960905097905906960512B90A98",
      INIT_12 => X"39068429704929999E999F9598598093559120990D3928090B60B9F81B990A49",
      INIT_13 => X"02A9A0439291D9099FC9C0044444450929790E90939D040491F90F90C029E002",
      INIT_14 => X"29290922C292CD20229F04392979081A2900202319104C2139F2824299204496",
      INIT_15 => X"09F009000940046F148005407096939F697692C64414469090097450343960C4",
      INIT_16 => X"8409930443403B9C7889288A23D88409A84A55A899EA9A85109E9B84109E9B84",
      INIT_17 => X"19E9C8A90E9C84A9E9D84CA9D89DA4E84D5A9E84C4E859810909F89410909F89",
      INIT_18 => X"4109099004C2590041901E9104419E91055190EE92059192E93892B293892294",
      INIT_19 => X"892B94045D829405950495095096059609960596054705197049709709804508",
      INIT_1A => X"09F8090809290C90C09019901990595A009A05A0459A09B059B09B09B0900000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
generic map (
      INIT_00 => X"D0A13102151E12E9EEF53E0EE1C40E8EE37771E1EE1A3E8EE141EFEEFB295FE0",
      INIT_01 => X"E229AFAFAFAF9EFA49E283E2EE3D44E16E142DE64F6EE16EC1DE61E6EE16E93D",
      INIT_02 => X"EACEE63DDEA5EEE687171EDE76DC18E144D1E666666419E83AE91AED5FE6EBE1",
      INIT_03 => X"CEE6FEE3E7081EE13333333CE91AE42DE6E5E5AE4CE85FE9E3E628FEE51AFF09",
      INIT_04 => X"DEFE345E7F3770E43E4A855E55EEE56E08A1E1BE74CCECDFE18E35BD2BEE13EB",
      INIT_05 => X"EEF1E317E0BBAEF2EF2EC71EBEFDEABE8EF61EBEFDE8BE6ED59E9A770EB7293E",
      INIT_06 => X"DE525E0E4470FD0E31E575EC2DE84E34E61ED5EA2E0571E33E5F4EC4EB310557",
      INIT_07 => X"91A5A69A01E9A1771EAA5EEDE072A59A4C56A19EFEDC9781757EFA5E23A5E5E1",
      INIT_08 => X"1E1E1E6FEEA5E553E06EB52A7EBE69E263E04EE45EEE56E19E52EAD66E13A0FD",
      INIT_09 => X"EFDC1193AE53A87E92ECA1E07EF3EF44A1E07E92F44D7E5145A46ECD7ED1EEE9",
      INIT_0A => X"72CBE3BFBE0C9E00E16E8E1C1E9EDB71EB0C56BE1BEE71E71A1EA1EE53EBA23B",
      INIT_0B => X"2810F2E755E09EFFDA0701E91E11E74491E11ED555FDE1655EFDED7A0E15DE5E",
      INIT_0C => X"E44AFBA19E85FE3E1F7B1B0C8DFE1EFF98AF81155E63E72DECE86EF06E86EE3E",
      INIT_0D => X"671EE40ED3E81E0F2FE9E565EDE8EA01EFD6F779A1E665811C52BE08A3E2252E",
      INIT_0E => X"A1EE62CA870AE55FED90E7EF620FA4295CE07C009EEE071E1D110933E09C1A32",
      INIT_0F => X"E84C9ECE915E9E344E0444560199FE1A5FF7E111D17E79D5BE08EE70E8E1775E",
      INIT_10 => X"E88EE3E2F5FDD17EE66CCF01379E9690E7A65EA3E6CE8A78AF68E188D5956E03",
      INIT_11 => X"E558EE07C0E1852D86EE1EE840E511B9D199EE23E6ADE4E9AE1FE840E56E8EE5",
      INIT_12 => X"2E891F5E75DE6EBDE8E8EFAFEEFEA3E018EF7DEE3B2E0A0E066DCEFC5CFE1EEE",
      INIT_13 => X"DCCE9542E6E54EDFEFBE625DDDDDDE5E1EAE12E5E2E6445EEA7710E5A11ED2A4",
      INIT_14 => X"3D2E5D41A3E2582A34EE442EAEFE7DF475179DA2BE667995BDF7A6F8E1D875E5",
      INIT_15 => X"6EE6DE3DDE3DAFF00FA86BA30DE2EFEF8E4AE1A8008DA1EAE1DE4D03090ED0AE",
      INIT_16 => X"A303ED4402A72CEDFDDEE5D4722B591E14E3DE63EE83EC4480E8E35980E8EB59",
      INIT_17 => X"8E8E323E08EB513E8E26558EA3E4310454E8E65CC1D62E751E7E22E651E7EC2E",
      INIT_18 => X"A51E7EE545990EF611ED58E68958E8EF8341E088E843E5E88E22E997EB1D32E2",
      INIT_19 => X"1E99E8954708EE44E673EA1EE1E12CE42CE82CEC4010429E45FE91ED3E061E13",
      INIT_1A => X"2EF82E1C2E00214111725EB38EF40DE32FE82EC5E8EF3E440E73EB3EE3E00000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000" )

